library ieee;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

--! 
package avalon_mem_pkg is
  
--	type t_mem_array is array(natural range <>) of std_logic_vector;

end package avalon_mem_pkg;
